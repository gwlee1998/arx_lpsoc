`ifndef __MUNOC_NODE_ID_H__
`define __MUNOC_NODE_ID_H__

`define NODE_ID_CORE_PERI_GROUP_NO_NAME (1)
`define NODE_ID_I_SNIM_I_SYSTEM_SRAM_NO_NAME (4)
`define NODE_ID_I_SNIM_COMMON_PERI_GROUP_NO_NAME (0)
`define NODE_ID_I_SNIM_EXTERNAL_PERI_GROUP_NO_NAME (2)
`define NODE_ID_I_SNIM_PLATFORM_CONTROLLER_NO_NAME (6)
`define NODE_ID_DEFAULT_SLAVE (15)
`define NODE_ID_I_MNIM_I_MAIN_CORE_INST (2)
`define NODE_ID_I_MNIM_I_MAIN_CORE_DATA_C (0)
`define NODE_ID_I_MNIM_I_MAIN_CORE_DATA_UC (1)
`define NODE_ID_I_MNIM_PLATFORM_CONTROLLER_MASTER (3)
`define NODE_ID_I_SNIM_I_USERIP1_SLAVE (5)
`define NODE_ID_I_SNIM_I_SYSTEM_DDR_NO_NAME (3)

`endif