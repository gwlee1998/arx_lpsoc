`ifndef __DCA_MODULE_MEMORYMAP_OFFSET_H__
`define __DCA_MODULE_MEMORYMAP_OFFSET_H__



// reg dca_matrix_lsu_inst_opcode
`define BW_DCA_MATRIX_LSU_INST_OPCODE 1
`define DCA_MATRIX_LSU_INST_OPCODE_DEFAULT_VALUE 0
`define DCA_MATRIX_LSU_INST_OPCODE_READ 0
`define DCA_MATRIX_LSU_INST_OPCODE_WRITE 1
`define DCA_MATRIX_LSU_INST_OPCODE_INDEX_WRITE 0

// reg dca_mru_inst
`define BW_DCA_MRU_INST 352
`define DCA_MRU_INST_DEFAULT_VALUE 0

// reg dca_mru_log
`define BW_DCA_MRU_LOG 32
`define DCA_MRU_LOG_DEFAULT_VALUE 0

// reg dca_mru_input
`define BW_DCA_MRU_INPUT 32
`define DCA_MRU_INPUT_DEFAULT_VALUE 0

// reg dca_mru_status
`define BW_DCA_MRU_STATUS 32
`define DCA_MRU_STATUS_DEFAULT_VALUE 0

// reg dca_mru_opcode
`define BW_DCA_MRU_OPCODE 5
`define DCA_MRU_OPCODE_DEFAULT_VALUE 0
`define DCA_MRU_OPCODE_NOP 1
`define DCA_MRU_OPCODE_COPY 2
`define DCA_MRU_OPCODE_TRANSPOSE 4
`define DCA_MRU_OPCODE_FILL 8
`define DCA_MRU_OPCODE_LSU0_REQ 16
`define DCA_MRU_OPCODE_INDEX_NOP 0
`define DCA_MRU_OPCODE_INDEX_COPY 1
`define DCA_MRU_OPCODE_INDEX_TRANSPOSE 2
`define DCA_MRU_OPCODE_INDEX_FILL 3
`define DCA_MRU_OPCODE_INDEX_LSU0_REQ 4
`define DCA_MRU_OPCODE_NONE 0

// reg dca_mru_fill_value
`define BW_DCA_MRU_FILL_VALUE 32
`define DCA_MRU_FILL_VALUE_DEFAULT_VALUE 0

// reg dca_matrix_mac_inst
`define BW_DCA_MATRIX_MAC_INST 512
`define DCA_MATRIX_MAC_INST_DEFAULT_VALUE 0

// reg dca_matrix_mac_log
`define BW_DCA_MATRIX_MAC_LOG 32
`define DCA_MATRIX_MAC_LOG_DEFAULT_VALUE 0

// reg dca_matrix_mac_status
`define BW_DCA_MATRIX_MAC_STATUS 32
`define DCA_MATRIX_MAC_STATUS_DEFAULT_VALUE 0

// reg dca_matrix_mac_opcode
`define BW_DCA_MATRIX_MAC_OPCODE 12
`define DCA_MATRIX_MAC_OPCODE_DEFAULT_VALUE 0
`define DCA_MATRIX_MAC_OPCODE_NO_CAL 1
`define DCA_MATRIX_MAC_OPCODE_ADDSUB 2
`define DCA_MATRIX_MAC_OPCODE_RSRC_INV 4
`define DCA_MATRIX_MAC_OPCODE_EWMULT 8
`define DCA_MATRIX_MAC_OPCODE_MULT_COND 16
`define DCA_MATRIX_MAC_OPCODE_INIT_ACC 32
`define DCA_MATRIX_MAC_OPCODE_LOAD_ACC 64
`define DCA_MATRIX_MAC_OPCODE_IS_FLOAT 128
`define DCA_MATRIX_MAC_OPCODE_LSU0_REQ 256
`define DCA_MATRIX_MAC_OPCODE_LSU1_REQ 512
`define DCA_MATRIX_MAC_OPCODE_LSU2_REQ 1024
`define DCA_MATRIX_MAC_OPCODE_RSRC_CONSTANT 2048
`define DCA_MATRIX_MAC_OPCODE_INDEX_NO_CAL 0
`define DCA_MATRIX_MAC_OPCODE_INDEX_ADDSUB 1
`define DCA_MATRIX_MAC_OPCODE_INDEX_RSRC_INV 2
`define DCA_MATRIX_MAC_OPCODE_INDEX_EWMULT 3
`define DCA_MATRIX_MAC_OPCODE_INDEX_MULT_COND 4
`define DCA_MATRIX_MAC_OPCODE_INDEX_INIT_ACC 5
`define DCA_MATRIX_MAC_OPCODE_INDEX_LOAD_ACC 6
`define DCA_MATRIX_MAC_OPCODE_INDEX_IS_FLOAT 7
`define DCA_MATRIX_MAC_OPCODE_INDEX_LSU0_REQ 8
`define DCA_MATRIX_MAC_OPCODE_INDEX_LSU1_REQ 9
`define DCA_MATRIX_MAC_OPCODE_INDEX_LSU2_REQ 10
`define DCA_MATRIX_MAC_OPCODE_INDEX_RSRC_CONSTANT 11
`define DCA_MATRIX_MAC_OPCODE_NONE 0

// reg dca_neugemm_inst
`define BW_DCA_NEUGEMM_INST 512
`define DCA_NEUGEMM_INST_DEFAULT_VALUE 0

// reg dca_neugemm_log
`define BW_DCA_NEUGEMM_LOG 32
`define DCA_NEUGEMM_LOG_DEFAULT_VALUE 0

// reg dca_neugemm_status
`define BW_DCA_NEUGEMM_STATUS 32
`define DCA_NEUGEMM_STATUS_DEFAULT_VALUE 0

// reg dca_neugemm_opcode
`define BW_DCA_NEUGEMM_OPCODE 13
`define DCA_NEUGEMM_OPCODE_DEFAULT_VALUE 0
`define DCA_NEUGEMM_OPCODE_NO_CAL 1
`define DCA_NEUGEMM_OPCODE_ADDSUB 2
`define DCA_NEUGEMM_OPCODE_RSRC_INV 4
`define DCA_NEUGEMM_OPCODE_EWMULT 8
`define DCA_NEUGEMM_OPCODE_MULT_COND 16
`define DCA_NEUGEMM_OPCODE_CONV_COND 32
`define DCA_NEUGEMM_OPCODE_INIT_ACC 64
`define DCA_NEUGEMM_OPCODE_LOAD_ACC 128
`define DCA_NEUGEMM_OPCODE_IS_FLOAT 256
`define DCA_NEUGEMM_OPCODE_LSU0_REQ 512
`define DCA_NEUGEMM_OPCODE_LSU1_REQ 1024
`define DCA_NEUGEMM_OPCODE_LSU2_REQ 2048
`define DCA_NEUGEMM_OPCODE_RSRC_CONSTANT 4096
`define DCA_NEUGEMM_OPCODE_INDEX_NO_CAL 0
`define DCA_NEUGEMM_OPCODE_INDEX_ADDSUB 1
`define DCA_NEUGEMM_OPCODE_INDEX_RSRC_INV 2
`define DCA_NEUGEMM_OPCODE_INDEX_EWMULT 3
`define DCA_NEUGEMM_OPCODE_INDEX_MULT_COND 4
`define DCA_NEUGEMM_OPCODE_INDEX_CONV_COND 5
`define DCA_NEUGEMM_OPCODE_INDEX_INIT_ACC 6
`define DCA_NEUGEMM_OPCODE_INDEX_LOAD_ACC 7
`define DCA_NEUGEMM_OPCODE_INDEX_IS_FLOAT 8
`define DCA_NEUGEMM_OPCODE_INDEX_LSU0_REQ 9
`define DCA_NEUGEMM_OPCODE_INDEX_LSU1_REQ 10
`define DCA_NEUGEMM_OPCODE_INDEX_LSU2_REQ 11
`define DCA_NEUGEMM_OPCODE_INDEX_RSRC_CONSTANT 12
`define DCA_NEUGEMM_OPCODE_NONE 0

// reg dca_neurgemm_inst
`define BW_DCA_NEURGEMM_INST 544
`define DCA_NEURGEMM_INST_DEFAULT_VALUE 0

// reg dca_neurgemm_log
`define BW_DCA_NEURGEMM_LOG 32
`define DCA_NEURGEMM_LOG_DEFAULT_VALUE 0

// reg dca_neurgemm_status
`define BW_DCA_NEURGEMM_STATUS 32
`define DCA_NEURGEMM_STATUS_DEFAULT_VALUE 0

// reg dca_neurgemm_opcode
`define BW_DCA_NEURGEMM_OPCODE 21
`define DCA_NEURGEMM_OPCODE_DEFAULT_VALUE 0
`define DCA_NEURGEMM_OPCODE_NO_CAL 1
`define DCA_NEURGEMM_OPCODE_ADDSUB 2
`define DCA_NEURGEMM_OPCODE_RSRC_INV 4
`define DCA_NEURGEMM_OPCODE_EWMULT 8
`define DCA_NEURGEMM_OPCODE_MULT_COND 16
`define DCA_NEURGEMM_OPCODE_CONV_COND 32
`define DCA_NEURGEMM_OPCODE_SEL_MAX 64
`define DCA_NEURGEMM_OPCODE_SEL_MIN 128
`define DCA_NEURGEMM_OPCODE_INIT_ACC 256
`define DCA_NEURGEMM_OPCODE_LOAD_ACC 512
`define DCA_NEURGEMM_OPCODE_IS_FLOAT 1024
`define DCA_NEURGEMM_OPCODE_LSU0_REQ 2048
`define DCA_NEURGEMM_OPCODE_LSU1_REQ 4096
`define DCA_NEURGEMM_OPCODE_LSU2_REQ 8192
`define DCA_NEURGEMM_OPCODE_RSRC_CONSTANT 16384
`define DCA_NEURGEMM_OPCODE_PAD_LOC_ROWU 32768
`define DCA_NEURGEMM_OPCODE_PAD_LOC_ROWD 65536
`define DCA_NEURGEMM_OPCODE_PAD_LOC_COLU 131072
`define DCA_NEURGEMM_OPCODE_PAD_LOC_COLD 262144
`define DCA_NEURGEMM_OPCODE_PAD_TYPE_ZERO 524288
`define DCA_NEURGEMM_OPCODE_OUTPUT_STRIDE 1048576
`define DCA_NEURGEMM_OPCODE_INDEX_NO_CAL 0
`define DCA_NEURGEMM_OPCODE_INDEX_ADDSUB 1
`define DCA_NEURGEMM_OPCODE_INDEX_RSRC_INV 2
`define DCA_NEURGEMM_OPCODE_INDEX_EWMULT 3
`define DCA_NEURGEMM_OPCODE_INDEX_MULT_COND 4
`define DCA_NEURGEMM_OPCODE_INDEX_CONV_COND 5
`define DCA_NEURGEMM_OPCODE_INDEX_SEL_MAX 6
`define DCA_NEURGEMM_OPCODE_INDEX_SEL_MIN 7
`define DCA_NEURGEMM_OPCODE_INDEX_INIT_ACC 8
`define DCA_NEURGEMM_OPCODE_INDEX_LOAD_ACC 9
`define DCA_NEURGEMM_OPCODE_INDEX_IS_FLOAT 10
`define DCA_NEURGEMM_OPCODE_INDEX_LSU0_REQ 11
`define DCA_NEURGEMM_OPCODE_INDEX_LSU1_REQ 12
`define DCA_NEURGEMM_OPCODE_INDEX_LSU2_REQ 13
`define DCA_NEURGEMM_OPCODE_INDEX_RSRC_CONSTANT 14
`define DCA_NEURGEMM_OPCODE_INDEX_PAD_LOC_ROWU 15
`define DCA_NEURGEMM_OPCODE_INDEX_PAD_LOC_ROWD 16
`define DCA_NEURGEMM_OPCODE_INDEX_PAD_LOC_COLU 17
`define DCA_NEURGEMM_OPCODE_INDEX_PAD_LOC_COLD 18
`define DCA_NEURGEMM_OPCODE_INDEX_PAD_TYPE_ZERO 19
`define DCA_NEURGEMM_OPCODE_INDEX_OUTPUT_STRIDE 20
`define DCA_NEURGEMM_OPCODE_NONE 0

`define BW_DCA_MATRIX_QDQ_INST 480
`define DCA_MATRIX_QDQ_INST_DEFAULT_VALUE 0

`define BW_DCA_MATRIX_QDQ_LOG 32
`define DCA_MATRIX_QDQ_LOG_DEFAULT_VALUE 0

`define BW_DCA_MATRIX_QDQ_STATUS 32
`define DCA_MATRIX_QDQ_STATUS_DEFAULT_VALUE 0

`endif
