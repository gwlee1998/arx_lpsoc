`ifndef __MUNOC_NODE_ID_H__
`define __MUNOC_NODE_ID_H__

`define NODE_ID_CORE_PERI_GROUP_NO_NAME (1)
`define NODE_ID_I_SNIM_I_SYSTEM_SRAM_NO_NAME (6)
`define NODE_ID_I_SNIM_COMMON_PERI_GROUP_NO_NAME (0)
`define NODE_ID_I_SNIM_EXTERNAL_PERI_GROUP_NO_NAME (2)
`define NODE_ID_I_SNIM_PLATFORM_CONTROLLER_NO_NAME (7)
`define NODE_ID_DEFAULT_SLAVE (15)
`define NODE_ID_I_SNIM_I_DCA_MATRIX_QGEMM_CONTROL_MMIOX1_INTERFACE_MMIO (4)
`define NODE_ID_I_MNIM_I_MAIN_CORE_INST (5)
`define NODE_ID_I_MNIM_I_MAIN_CORE_DATA_C (3)
`define NODE_ID_I_MNIM_I_MAIN_CORE_DATA_UC (4)
`define NODE_ID_I_MNIM_PLATFORM_CONTROLLER_MASTER (6)
`define NODE_ID_I_MNIM_I_DCA_MATRIX_QGEMM_MX_MLSU_NOC_PART (2)
`define NODE_ID_I_MNIM_I_DCA_MATRIX_QGEMM_MW_MLSU_NOC_PART (1)
`define NODE_ID_I_MNIM_I_DCA_MATRIX_QGEMM_MO_MLSU_NOC_PART (0)
`define NODE_ID_I_SNIM_I_DCA_MATRIX_QGEMM_MQ2VTA (3)
`define NODE_ID_I_SNIM_I_SYSTEM_DDR_NO_NAME (5)

`endif