`ifndef __MEMORYMAP_INFO_H__
`define __MEMORYMAP_INFO_H__


`define I_SYSTEM_DDR_BASEADDR (32'h 0)
`define I_SYSTEM_DDR_SIZE (32'h 40000000)
`define I_SYSTEM_DDR_LASTADDR (32'h 3fffffff)
`define I_USERIP1_SLAVE_BASEADDR (32'h c0000000)
`define I_USERIP1_SLAVE_SIZE (32'h 8000)
`define I_USERIP1_SLAVE_LASTADDR (32'h c0007fff)
`define DEFAULT_SLAVE_BASEADDR (32'h c0008000)
`define DEFAULT_SLAVE_SIZE (32'h 1000)
`define DEFAULT_SLAVE_LASTADDR (32'h c0008fff)
`define I_SYSTEM_SRAM_BASEADDR (32'h e0000000)
`define I_SYSTEM_SRAM_SIZE (32'h 8000)
`define I_SYSTEM_SRAM_LASTADDR (32'h e0007fff)
`define PLATFORM_CONTROLLER_BASEADDR (32'h e1000000)
`define PLATFORM_CONTROLLER_SIZE (32'h 40000)
`define PLATFORM_CONTROLLER_LASTADDR (32'h e103ffff)
`define COMMON_PERI_GROUP_BASEADDR (32'h e2000000)
`define COMMON_PERI_GROUP_SIZE (32'h 10000)
`define COMMON_PERI_GROUP_LASTADDR (32'h e200ffff)
`define EXTERNAL_PERI_GROUP_BASEADDR (32'h e2010000)
`define EXTERNAL_PERI_GROUP_SIZE (32'h 10000)
`define EXTERNAL_PERI_GROUP_LASTADDR (32'h e201ffff)
`define CORE_PERI_GROUP_BASEADDR (32'h f0000000)
`define CORE_PERI_GROUP_SIZE (32'h 8000)
`define CORE_PERI_GROUP_LASTADDR (32'h f0007fff)
`define NOC_CONTROLLER_BASEADDR (32'h c0008000)
`define IROM_BASEADDR (32'h e2000000)

`endif