case(NETWORK_TYPE)
	`FORWARD_NETWORK:
		case(ROUTER_ID)
			`ROUTER_ID_I_SYSTEM_ROUTER:
				case(target_node)
					`NODE_ID_I_SNIM_I_SYSTEM_SRAM_NO_NAME: routing_info = 6'b 000001;
					`NODE_ID_I_SNIM_COMMON_PERI_GROUP_NO_NAME: routing_info = 6'b 000010;
					`NODE_ID_I_SNIM_EXTERNAL_PERI_GROUP_NO_NAME: routing_info = 6'b 000100;
					`NODE_ID_I_SNIM_PLATFORM_CONTROLLER_NO_NAME: routing_info = 6'b 001000;
					`NODE_ID_DEFAULT_SLAVE: routing_info = 6'b 010000;
					`NODE_ID_I_SNIM_I_DCA_MATRIX_QGEMM_CONTROL_MMIOX1_INTERFACE_MMIO: routing_info = 6'b 100000;
				endcase
			`ROUTER_ID_I_USER_ROUTER:
				case(target_node)
					`NODE_ID_I_SNIM_I_DCA_MATRIX_QGEMM_MQ2VTA: routing_info = 8'b 00000001;
					`NODE_ID_I_SNIM_I_SYSTEM_DDR_NO_NAME: routing_info = 8'b 00000010;
					`NODE_ID_I_SNIM_I_SYSTEM_SRAM_NO_NAME: routing_info = 8'b 00000100;
					`NODE_ID_I_SNIM_COMMON_PERI_GROUP_NO_NAME: routing_info = 8'b 00000100;
					`NODE_ID_I_SNIM_EXTERNAL_PERI_GROUP_NO_NAME: routing_info = 8'b 00000100;
					`NODE_ID_I_SNIM_PLATFORM_CONTROLLER_NO_NAME: routing_info = 8'b 00000100;
					`NODE_ID_DEFAULT_SLAVE: routing_info = 8'b 00000100;
					`NODE_ID_I_SNIM_I_DCA_MATRIX_QGEMM_CONTROL_MMIOX1_INTERFACE_MMIO: routing_info = 8'b 00000100;
				endcase
		endcase
	`BACKWARD_NETWORK:
		case(ROUTER_ID)
			`ROUTER_ID_I_SYSTEM_ROUTER:
				case(target_node)
					`NODE_ID_I_MNIM_I_MAIN_CORE_INST: routing_info = 7'b 0000001;
					`NODE_ID_I_MNIM_I_MAIN_CORE_DATA_C: routing_info = 7'b 0000001;
					`NODE_ID_I_MNIM_I_MAIN_CORE_DATA_UC: routing_info = 7'b 0000001;
					`NODE_ID_I_MNIM_PLATFORM_CONTROLLER_MASTER: routing_info = 7'b 0000001;
					`NODE_ID_I_MNIM_I_DCA_MATRIX_QGEMM_MX_MLSU_NOC_PART: routing_info = 7'b 0000001;
					`NODE_ID_I_MNIM_I_DCA_MATRIX_QGEMM_MW_MLSU_NOC_PART: routing_info = 7'b 0000001;
					`NODE_ID_I_MNIM_I_DCA_MATRIX_QGEMM_MO_MLSU_NOC_PART: routing_info = 7'b 0000001;
				endcase
			`ROUTER_ID_I_USER_ROUTER:
				case(target_node)
					`NODE_ID_I_MNIM_I_MAIN_CORE_INST: routing_info = 7'b 0000001;
					`NODE_ID_I_MNIM_I_MAIN_CORE_DATA_C: routing_info = 7'b 0000010;
					`NODE_ID_I_MNIM_I_MAIN_CORE_DATA_UC: routing_info = 7'b 0000100;
					`NODE_ID_I_MNIM_PLATFORM_CONTROLLER_MASTER: routing_info = 7'b 0001000;
					`NODE_ID_I_MNIM_I_DCA_MATRIX_QGEMM_MX_MLSU_NOC_PART: routing_info = 7'b 0010000;
					`NODE_ID_I_MNIM_I_DCA_MATRIX_QGEMM_MW_MLSU_NOC_PART: routing_info = 7'b 0100000;
					`NODE_ID_I_MNIM_I_DCA_MATRIX_QGEMM_MO_MLSU_NOC_PART: routing_info = 7'b 1000000;
				endcase
		endcase
endcase